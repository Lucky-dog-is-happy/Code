module connect(
	input wire sw,
	output wire led
);
	assign led = sw;
endmodule